H2O                                     
   1.00000000000000     
    -8.0330016028837967    8.0329698381748678    8.0329698602708426
     8.0329698602708390   -8.0330016028837985    8.0329698381748660
     8.0329698381748660    8.0329698602708426   -8.0330016028837985
   H    O 
    96    48
Direct
  0.9478240946061267  0.2225293515463579  0.0717545105210136
  0.6239268560808297  0.2747018783133879  0.5521825880428397
  0.6507759405780441  0.8760764226513761  0.4282580787469047
  0.2747018783133879  0.5521825880428397  0.6239268560808297
  0.7252987178160072  0.7774788161602255  0.3492212895737077
  0.4478238141000036  0.5717526162013570  0.7225263499884998
  0.9478182153652677  0.2252929156083347  0.8760785665885494
  0.7747022470739783  0.1507714055770335  0.7225253734668957
  0.4282506164642325  0.2774789647290439  0.5521785206380394
  0.6507734999423088  0.2746992318588272  0.2225220218729218
  0.4282580787469047  0.6507759405780441  0.8760764226513761
  0.7225253734668957  0.7747022470739783  0.1507714055770335
  0.1507714055770335  0.7225253734668957  0.7747022470739783
  0.9282562291798898  0.0521805100533727  0.7774809723986842
  0.8492321755430303  0.0717529153255767  0.6239325486057258
  0.0521805100533727  0.7774809723986842  0.9282562291798898
  0.2746992318588272  0.2225220218729218  0.6507734999423088
  0.0717545105203599  0.9478240946057928  0.2225293515460808
  0.0521801012414401  0.7746979482559526  0.1239302173768911
  0.2225220218729218  0.6507734999423088  0.2746992318588272
  0.7225263499884998  0.4478238141000036  0.5717526162013570
  0.4478231945396405  0.3760704233363308  0.7252954061696970
  0.6239325486057258  0.8492321755430303  0.0717529153255767
  0.9282496753151012  0.3760743465909127  0.1507831622441751
  0.3760704233363308  0.7252954061696970  0.4478231945396405
  0.1239216749768878  0.5717394468959758  0.3492159641588543
  0.2253008329966352  0.8492226940536793  0.2774770098768003
  0.8760764226513761  0.4282580787469047  0.6507759405780441
  0.5521785206380394  0.4282506164642325  0.2774789647290439
  0.2774770098768003  0.2253008329966352  0.8492226940536793
  0.7252954061696970  0.4478231945396405  0.3760704233363308
  0.8760785665885494  0.9478182153652677  0.2252929156083347
  0.3760743465909127  0.1507831622441751  0.9282496753151012
  0.3492159641588543  0.1239216749768878  0.5717394468959758
  0.7774809723986842  0.9282562291798898  0.0521805100533727
  0.7746979482559526  0.1239302173768911  0.0521801012414401
  0.1507831622441751  0.9282496753151012  0.3760743465909127
  0.0717529153255767  0.6239325486057258  0.8492321755430303
  0.1239302173768911  0.0521801012414401  0.7746979482559526
  0.2774789647290439  0.5521785206380394  0.4282506164642325
  0.3492212895737077  0.7252987178160072  0.7774788161602255
  0.2225293515460808  0.0717545105203599  0.9478240946057928
  0.7774788161602255  0.3492212895737077  0.7252987178160072
  0.5521825880428397  0.6239268560808297  0.2747018783133879
  0.8492226940536793  0.2774770098768003  0.2253008329966352
  0.2252929156083347  0.8760785665885494  0.9478182153652677
  0.5717394468959758  0.3492159641588543  0.1239216749768878
  0.5717526162013570  0.7225263499884998  0.4478238141000036
  0.9130453794822458  0.1085208988393675  0.9645823929922993
  0.5515297948100041  0.1954751067327665  0.5869600367990734
  0.6439484997152055  0.9484719583780422  0.5354364556003072
  0.1954751067327665  0.5869600367990734  0.5515297948100041
  0.8045230403608032  0.8914859842414833  0.3560555573350184
  0.4130385124498563  0.4645746456618649  0.6085160528432026
  0.9130353316832357  0.3045210840723837  0.9484700706919679
  0.6954730756383657  0.1439381506146150  0.6085172909400270
  0.5354290852731837  0.3914855331792256  0.5869603884468957
  0.6439424023385676  0.1954739009176185  0.1085185365914030
  0.5354364556003072  0.6439484997152055  0.9484719583780422
  0.6085172909400270  0.6954730756383657  0.1439381506146150
  0.1439381506146150  0.6085172909400270  0.6954730756383657
  0.0354313508361228  0.0869652086629100  0.8914882861766875
  0.8560607191268800  0.9645777535396945  0.5515348591181913
  0.0869652086629100  0.8914882861766875  0.0354313508361228
  0.1954739009176185  0.1085185365914030  0.6439424023385676
  0.9645823929921856  0.9130453794821748  0.1085208988393888
  0.0869623402079165  0.6954742896506937  0.0515354092403432
  0.1085185365914030  0.6439424023385676  0.1954739009176185
  0.6085160528432026  0.4130385124498563  0.4645746456618649
  0.4130437553472410  0.4484685238382817  0.8045224707710970
  0.5515348591181913  0.8560607191268800  0.9645777535396945
  0.0354209858716816  0.4484665003056242  0.1439423365106106
  0.4484685238382817  0.8045224707710970  0.4130437553472410
  0.0515314198485353  0.4645663667475685  0.3560545730794166
  0.3045267382536376  0.8560571128219517  0.3914854428280840
  0.9484719583780422  0.5354364556003072  0.6439484997152055
  0.5869603884468957  0.5354290852731837  0.3914855331792256
  0.3914854428280840  0.3045267382536376  0.8560571128219517
  0.8045224707710970  0.4130437553472410  0.4484685238382817
  0.9484700706919679  0.9130353316832357  0.3045210840723837
  0.4484665003056242  0.1439423365106106  0.0354209858716816
  0.3560545730794166  0.0515314198485353  0.4645663667475685
  0.8914882861766875  0.0354313508361228  0.0869652086629100
  0.6954742896506937  0.0515354092403432  0.0869623402079165
  0.1439423365106106  0.0354209858716816  0.4484665003056242
  0.9645777535396945  0.5515348591181913  0.8560607191268800
  0.0515354092403432  0.0869623402079165  0.6954742896506937
  0.3914855331792256  0.5869603884468957  0.5354290852731837
  0.3560555573350184  0.8045230403608032  0.8914859842414833
  0.1085208988393888  0.9645823929921856  0.9130453794821748
  0.8914859842414833  0.3560555573350184  0.8045230403608032
  0.5869600367990734  0.5515297948100041  0.1954751067327665
  0.8560571128219517  0.3914854428280840  0.3045267382536376
  0.3045210840723837  0.9484700706919679  0.9130353316832357
  0.4645663667475685  0.3560545730794166  0.0515314198485353
  0.4645746456618649  0.6085160528432026  0.4130385124498563
  0.9049749384637863  0.1370631592265569  0.0342433066535540
  0.6292663997712922  0.2320988133752248  0.5950455709940637
  0.6028316548863065  0.8707375868428590  0.4657796581778776
  0.2320988133752248  0.5950455709940637  0.6292663997712922
  0.7679057833994611  0.8629447809086763  0.3971710351313559
  0.4049635821991072  0.5342320359464514  0.6370601681535218
  0.9049584783350892  0.2678992799408969  0.8707369273967938
  0.7320950697141787  0.1028259789682111  0.6370588491131005
  0.4657739559769222  0.3629453265133402  0.5950399398660039
  0.6028281459537537  0.2320960236111855  0.1370561782318452
  0.4657796581778776  0.6028316548863065  0.8707375868428590
  0.6370588491131005  0.7320950697141787  0.1028259789682111
  0.1028259789682111  0.6370588491131005  0.7320950697141787
  0.9657782693559074  0.0950471590430058  0.8629468330127159
  0.8971786585034044  0.0342337293754859  0.6292693969696503
  0.0950471590430058  0.8629468330127159  0.9657782693559074
  0.2320960236111855  0.1370561782318452  0.6028281459537537
  0.0342433066541580  0.9049749384640847  0.1370631592268553
  0.0950353276438764  0.7320878169500639  0.1292682168745407
  0.1370561782318452  0.6028281459537537  0.2320960236111855
  0.6370601681535218  0.4049635821991072  0.5342320359464514
  0.4049643381281203  0.3707338999269499  0.7679027079252242
  0.6292693969696503  0.8971786585034044  0.0342337293754859
  0.9657644971541380  0.3707335866953775  0.1028317968135914
  0.3707338999269499  0.7679027079252242  0.4049643381281203
  0.1292635799489327  0.5342243464123749  0.3971664450635706
  0.2679093216611899  0.8971727055993919  0.3629427949238282
  0.8707375868428590  0.4657796581778776  0.6028316548863065
  0.5950399398660039  0.4657739559769222  0.3629453265133402
  0.3629427949238282  0.2679093216611899  0.8971727055993919
  0.7679027079252242  0.4049643381281203  0.3707338999269499
  0.8707369273967938  0.9049584783350892  0.2678992799408969
  0.3707335866953775  0.1028317968135914  0.9657644971541380
  0.3971664450635706  0.1292635799489327  0.5342243464123749
  0.8629468330127159  0.9657782693559074  0.0950471590430058
  0.7320878169500639  0.1292682168745407  0.0950353276438764
  0.1028317968135914  0.9657644971541380  0.3707335866953775
  0.0342337293754859  0.6292693969696503  0.8971786585034044
  0.1292682168745407  0.0950353276438764  0.7320878169500639
  0.3629453265133402  0.5950399398660039  0.4657739559769222
  0.3971710351313559  0.7679057833994611  0.8629447809086763
  0.1370631592268553  0.0342433066541580  0.9049749384640847
  0.8629447809086763  0.3971710351313559  0.7679057833994611
  0.5950455709940637  0.6292663997712922  0.2320988133752248
  0.8971727055993919  0.3629427949238282  0.2679093216611899
  0.2678992799408969  0.8707369273967938  0.9049584783350892
  0.5342243464123749  0.3971664450635706  0.1292635799489327
  0.5342320359464514  0.6370601681535218  0.4049635821991072
 
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
  0.00000000E+00  0.00000000E+00  0.00000000E+00
